LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MUX2_1 IS
	PORT(A, B, SEL : IN STD_LOGIC;
				F,C : OUT STD_LOGIC);
END MUX2_1;

ARCHITECTURE BEHAVIORAL OF MUX2_1 IS

BEGIN
	WITH SEL SELECT
		F<=A WHEN '0',
			B WHEN '1',
			'0' WHEN OTHERS;
END BEHAVIORAL;