LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MUX10TO1 IS
	PORT(R0: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			R1: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			R2: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			R3: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			R4: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			R5: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			R6: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			R7: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			DIN: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			GIN: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			SEL: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			Q: OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
END MUX10TO1;

ARCHITECTURE BEHAVIORAL OF MUX10TO1 IS
	BEGIN
		PROCESS(SEL,R0,R1,R2,R3,R4,R5,R6,R7,DIN,GIN)
		BEGIN
			CASE SEL IS
				WHEN "0000" =>
					Q<=R0;
				WHEN "0001" =>
					Q<=R1;
				WHEN "0010" =>
					Q<=R2;
				WHEN "0011" =>
					Q<=R3;
				WHEN "0100" =>
					Q<=R4;
				WHEN "0101" =>
					Q<=R5;
				WHEN "0110" =>
					Q<=R6;
				WHEN "0111" =>
					Q<=R7;
				WHEN "1000" =>
					Q<=DIN;
				WHEN "1001" =>
					Q<=GIN;
				WHEN OTHERS =>
					Q<="000000000";
			END CASE;
		END PROCESS;
END BEHAVIORAL;
			