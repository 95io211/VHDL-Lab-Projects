LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ENCODER IS
	PORT(A: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
			Q: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENCODER;

ARCHITECTURE BEHAVIORAL OF ENCODER IS
BEGIN
	PROCESS(A)
	BEGIN
		CASE A IS 
			WHEN "0000000001" => Q<="0000";
			WHEN "0000000010" => Q<="0001";
			WHEN "0000000100" => Q<="0010";
			WHEN "0000001000" => Q<="0011";
			WHEN "0000010000" => Q<="0100";
			WHEN "0000100000" => Q<="0101";
			WHEN "0001000000" => Q<="0110";
			WHEN "0010000000" => Q<="0111";
			WHEN "0100000000" => Q<="1000";
			WHEN "1000000000" => Q<="1001";
			WHEN OTHERS => Q <="0000";
		END CASE;
	END PROCESS;
END BEHAVIORAL;