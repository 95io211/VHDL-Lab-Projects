LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY BEHAVIORALDIVIDER IS
	PORT(DIVIDEND: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			DIVISOR: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			QUOTIENT: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			REMAINDER: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END BEHAVIORALDIVIDER;

ARCHITECTURE BEHAVIORAL OF BEHAVIORALDIVIDER IS

BEGIN
PROCESS(DIVIDEND,DIVISOR)
VARIABLE COUNTER: STD_LOGIC_VECTOR(9 DOWNTO 0);
VARIABLE REMAINS: STD_LOGIC_VECTOR(15 DOWNTO 0);
BEGIN
	IF DIVIDEND = DIVISOR THEN
		REMAINS:=(OTHERS=>'0');
		COUNTER:="0000000001";
	ELSIF DIVIDEND < DIVISOR THEN
		REMAINS:=DIVIDEND;
		COUNTER:="0000000000";
	ELSIF DIVIDEND > DIVISOR THEN
	REMAINS:=DIVIDEND;
	COUNTER:="0000000000";
		WHILE ((REMAINS >= DIVISOR) AND COUNTER<"1111111111") LOOP
			REMAINS:=REMAINS-DIVISOR;
			COUNTER:=COUNTER+"0000000001";
		END LOOP;
	END IF;
REMAINDER<=REMAINS;
QUOTIENT<=COUNTER;
END PROCESS;
END BEHAVIORAL;