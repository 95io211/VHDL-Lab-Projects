LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY DECODER IS
	PORT(A: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			Q: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END DECODER;

ARCHITECTURE BEHAVIORAL OF DECODER IS
BEGIN
	PROCESS(A)
	BEGIN
		CASE A IS 
			WHEN "000" => Q<="00000001";
			WHEN "001" => Q<="00000010";
			WHEN "010" => Q<="00000100";
			WHEN "011" => Q<="00001000";
			WHEN "100" => Q<="00010000";
			WHEN "101" => Q<="00100000";
			WHEN "110" => Q<="01000000";
			WHEN "111" => Q<="10000000";
			WHEN OTHERS => Q <="00000000";
		END CASE;
	END PROCESS;
END BEHAVIORAL;