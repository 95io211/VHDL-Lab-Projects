LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY REGISTERS8 IS
	PORT(DR0: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			DR1: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			DR2: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			DR3: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			DR4: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			DR5: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			DR6: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			DR7: IN STD_LOGIC_VECTOR(8 DOWNTO 0);
			clk,R0,R1,R2,R3,R4,R5,R6,R7,R8: IN STD_LOGIC;
			OR0: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
			OR1: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
			OR2: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
			OR3: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
			OR4: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
			OR5: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
			OR6: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
			OR7: OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
END REGISTERS8;

ARCHITECTURE BEHAVIORAL OF REGISTERS8 IS

BEGIN
	PROCESS(clk,R1,R2,R3,R4,R5,R6,R7,DR1,DR2,DR3,DR4,DR5,DR6,DR7)
	BEGIN
		IF clk'EVENT AND clk='1' THEN
			IF R0='1' THEN
				OR0<=DR0;
			ELSIF R1='1' THEN
				OR1<=DR1;
			ELSIF R2='1' THEN
				OR2<=DR2;
			ELSIF R3='1' THEN
				OR3<=DR3;
			ELSIF R4='1' THEN
				OR4<=DR4;
			ELSIF R5='1' THEN
				OR5<=DR5;
			ELSIF R6='1' THEN
				OR6<=DR6;
			ELSIF R7='1' THEN
				OR7<=DR7;
			END IF;
		END IF;
	END PROCESS;
END BEHAVIORAL;