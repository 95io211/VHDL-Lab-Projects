LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ROM64x16 IS
	PORT(ADDRESS: IN INTEGER RANGE 0 TO 7;
			DATA: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END ROM64x16;

ARCHITECTURE BEHAVIORAL OF ROM64x16 IS
	TYPE ROM_ARRAY IS ARRAY(0 TO 7) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	CONSTANT ROM: ROM_ARRAY:=( "00000",
										"00001",
										"00010",
										"00011",
										"00100",
										"00101",
										"00110",
										"00111");
	
	BEGIN
		DATA<=ROM(ADDRESS);
END BEHAVIORAL;